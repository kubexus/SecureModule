----------------------------------
-- Łukasz DZIEŁ (883533374)     --
-- FPGACOMMEXAMPLE-v2           --
-- 01.2016                      --
-- 1.0                          --
----------------------------------

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY RS232_STANDARD_INTERFACE IS PORT
(	
	CLK	:IN STD_LOGIC;
	INIT	:IN STD_LOGIC;
	
	TX		:OUT STD_LOGIC;
	RX		:IN STD_LOGIC;
	
	INT_WR		:OUT STD_LOGIC;
	INT_RD		:OUT STD_LOGIC;
	INT_ADDR		:OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
	INT_DIN		:IN STD_LOGIC_VECTOR(31 DOWNTO 0);
	INT_DOUT		:OUT STD_LOGIC_VECTOR(31 DOWNTO 0)
);
END ENTITY;

ARCHITECTURE RS232_STANDARD_INTERFACE_ARCH OF RS232_STANDARD_INTERFACE IS
	
	SIGNAL TEMP0 :STD_LOGIC;
	SIGNAL TEMP1 :STD_LOGIC;
	SIGNAL TEMP2 :STD_LOGIC;
	SIGNAL TEMP3 :STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL TEMP4 :STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN
	unit01 : ENTITY WORK.RS232_INTERFACE PORT MAP (CLK, INIT, TX, TEMP0, TEMP4, RX, TEMP1, TEMP2, TEMP3);
	unit02 : ENTITY WORK.COMMAND_CONTROL PORT MAP (CLK, INIT, TEMP2, TEMP1, TEMP0, TEMP3, TEMP4,
																	INT_WR, INT_RD, INT_ADDR, INT_DIN, INT_DOUT);
END ARCHITECTURE;